module m21(D0, D1, S, Y);
	output Y;
	input D0, D1, S;

	assign Y=S?D1:D0;

endmodule
